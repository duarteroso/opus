module file

#flag linux -I/usr/include/opus
#flag linux -lopusfile

#include "opusfile.h"
