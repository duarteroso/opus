module file

pub const op_false = -1
pub const op_eof = -2
pub const op_hole = -3
pub const op_eread = -128
pub const op_efault = -129
pub const op_eimpl = -130
pub const op_einval = -131
pub const op_enotformat = -132
pub const op_ebadheader = -133
pub const op_eversion = -134
pub const op_enotaudio = -135
pub const op_ebadpacket = -136
pub const op_ebadlink = -137
pub const op_enoseek = -138
pub const op_ebadtimestamp = -139
pub const opus_channel_count_max = 255

pub const chunk = 4096
