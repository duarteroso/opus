module file

#flag linux -lopusfile

#flag darwin -I/usr/local/opt/opusfile/include/opus
#flag darwin -I/usr/local/opt/opus/include/opus
#flag darwin -L/usr/local/opt/opusfile/lib
#flag darwin -lopusfile

#include "opusfile.h"
